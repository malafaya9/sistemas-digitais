library verilog;
use verilog.vl_types.all;
entity REG16_vlg_vec_tst is
end REG16_vlg_vec_tst;
