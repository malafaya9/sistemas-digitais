library verilog;
use verilog.vl_types.all;
entity ADD1_vlg_vec_tst is
end ADD1_vlg_vec_tst;
