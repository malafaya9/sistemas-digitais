library verilog;
use verilog.vl_types.all;
entity CTL2000_vlg_vec_tst is
end CTL2000_vlg_vec_tst;
