library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Controlador is 
	port
	(
	clk:in std_logic
	);
end Controlador;
architecture behavioral of Controlador is
begin
	process(clk)
	begin
		
	end process;
end behavioral;