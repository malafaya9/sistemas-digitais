library verilog;
use verilog.vl_types.all;
entity MUX5E_vlg_vec_tst is
end MUX5E_vlg_vec_tst;
