library verilog;
use verilog.vl_types.all;
entity COMP_vlg_vec_tst is
end COMP_vlg_vec_tst;
