library verilog;
use verilog.vl_types.all;
entity COMP0_vlg_check_tst is
    port(
        out_comp        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end COMP0_vlg_check_tst;
