library ieee;
use ieee.std_logic_1164.all;

entity MUX4E is
  port(
    sel : in std_logic_vector(1 downto 0);                      
    a   : in std_logic_vector(7 downto 0);   
    b   : in std_logic_vector(7 downto 0);
	 c   : in std_logic_vector(7 downto 0);
	 d   : in std_logic_vector(7 downto 0);
	 --y   : in std_logic_vector(9 downto 0);	 
	 out_mux : out std_logic_vector(7 downto 0) 
    
  );
end MUX4E;


architecture dataflow of MUX4E is

begin
  process(sel, a, b, c, d)
  begin
	case sel is
		when "00" =>
			out_mux <= a;
		when "01" =>
			out_mux <= b;
		when "10" =>
			out_mux <= c;
		when "11" =>
			out_mux <= d;
	end case;
  end process;

end dataflow;