library verilog;
use verilog.vl_types.all;
entity MUX2E_vlg_vec_tst is
end MUX2E_vlg_vec_tst;
