library verilog;
use verilog.vl_types.all;
entity MEMDATA_vlg_vec_tst is
end MEMDATA_vlg_vec_tst;
