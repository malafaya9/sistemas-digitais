library verilog;
use verilog.vl_types.all;
entity COMP0_vlg_vec_tst is
end COMP0_vlg_vec_tst;
