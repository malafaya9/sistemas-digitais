library verilog;
use verilog.vl_types.all;
entity REG8_vlg_vec_tst is
end REG8_vlg_vec_tst;
