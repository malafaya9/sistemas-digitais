library verilog;
use verilog.vl_types.all;
entity MUX4E_vlg_vec_tst is
end MUX4E_vlg_vec_tst;
